module M();

    initial
    accept_on
        begin
            11_11
            -11_11
            12'sb0101101
