module M();

    initial
        begin
            $display("Hello World");
        end

endmodule
